module xor_gate (
input a,b,
output y);

   xor x1(y,a,b); 
endmodule
